video_PLL_inst : video_PLL PORT MAP (
		inclk0	 => inclk0_sig,
		c0	 => c0_sig
	);
