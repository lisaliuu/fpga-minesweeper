LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

Entity board is (
	Port (

	)
)

-- Board is a 8x8 grid of squares
-- 01 02 03 04 05 06 07 08
-- 09 10 11 12 13 14 15 16
-- 17 18 19 20 21 22 23 24
-- 25 26 27 28 29 30 31 32
-- 33 34 35 36 37 38 39 40
-- 41 42 43 44 45 46 47 48
-- 49 50 51 52 53 54 55 56
-- 57 58 59 60 61 62 63 64