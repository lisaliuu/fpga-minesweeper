LIBRARY ieee;
USE ieee.std_logic_1164.ALL;

ENTITY bcd_seven IS
	PORT
	(
		bcd : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		H0 : OUT STD_LOGIC_VECTOR(6 DOWNTO 0)
	);
END bcd_seven;

ARCHITECTURE behavioral OF bcd_seven IS
BEGIN
	WITH bcd SELECT H0 <=
		"1000000" WHEN "0000",
		"1111001" WHEN "0001",
		"0100100" WHEN "0010",
		"0110000" WHEN "0011",
		"0011001" WHEN "0100",
		"0010010" WHEN "0101",
		"0000010" WHEN "0110",
		"1111000" WHEN "0111",
		"0000000" WHEN "1000",
		"0010000" WHEN "1001",
		"0111111" WHEN OTHERS;
END behavioral;