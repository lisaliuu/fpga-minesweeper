LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

USE work.board_layout_pkg.ALL;

ENTITY board IS
	PORT
	(
		Vert_sync, Horiz_sync : IN STD_LOGIC;
		pixel_row, pixel_column : IN STD_LOGIC_VECTOR(9 DOWNTO 0);
		Red, Green, Blue : OUT STD_LOGIC;
		-- signals from logic
		cell_status : IN board_bool;
		cell_flagged : IN board_bool;
		cell_value : IN board_size;
		cell_userb : IN user_pos
	);
END board;

-- Board is a 8x8 grid of squares
-- 50 x 50 pixels for each square
-- 640 x 480 (WIDTH = 640, HEIGHT = 480)
-- |                   four pixels                 |
-- | <= 84 => | 01 02 03 04 05 06 07 08 | <= 84 => | 00 01 02 03 04 05 06 07
-- | <= 84 => | 09 10 11 12 13 14 15 16 | <= 84 => | 10 11 12 13 14 15 16 17
-- | <= 84 => | 17 18 19 20 21 22 23 24 | <= 84 => | 20 21 22 23 24 25 26 27
-- | <= 84 => | 25 26 27 28 29 30 31 32 | <= 84 => | 30 31 32 33 34 35 36 37
-- | <= 84 => | 33 34 35 36 37 38 39 40 | <= 84 => | 40 41 42 43 44 45 46 47
-- | <= 84 => | 41 42 43 44 45 46 47 48 | <= 84 => | 50 51 52 53 54 55 56 57
-- | <= 84 => | 49 50 51 52 53 54 55 56 | <= 84 => | 60 61 62 63 64 65 66 67
-- | <= 84 => | 57 58 59 60 61 62 63 64 | <= 84 => | 70 71 72 73 74 75 76 77
-- |                   four pixels                 |

-- w = h = 50
-- 0-83 || 84-91 | "92-141", 142-149, "150-199", 200-207, "208-257", 258-265, "266-315", 316-323, "324-373", 374-381, "382-431", 432-439, "440-489", 490-497, "498-547" | 548-555 || 556-639
-- e.g.  01 (91,  4) < (x, y) < (142,  4) | 02 (140) ...
--          (91, 54) < (x, y) < (142, 54) |    (140) ...
ARCHITECTURE behavior OF board IS
	-- Video Display Signals
	--MARK: signal for colors
	SIGNAL background_color : STD_LOGIC_VECTOR(2 DOWNTO 0) := "111"; -- white
	SIGNAL grid_color : STD_LOGIC_VECTOR(2 DOWNTO 0) := "000"; -- black
	SIGNAL opened_cell_color : STD_LOGIC_VECTOR(2 DOWNTO 0) := "000"; -- black
	SIGNAL closed_cell_color : STD_LOGIC_VECTOR(2 DOWNTO 0) := "010"; -- green
	SIGNAL flagged_cell_color : STD_LOGIC_VECTOR(2 DOWNTO 0) := "100"; -- red
	--MARK: signal for display
	SIGNAL display_width : STD_LOGIC_VECTOR(9 DOWNTO 0) := CONV_STD_LOGIC_VECTOR(640, 10);
	SIGNAL display_height : STD_LOGIC_VECTOR(9 DOWNTO 0) := CONV_STD_LOGIC_VECTOR(480, 10);
	--MARK: signal for background
	SIGNAL margin_width, margin_height : STD_LOGIC_VECTOR(9 DOWNTO 0) := CONV_STD_LOGIC_VECTOR(472, 10); -- 50*8+8*9
	SIGNAL margin_x : STD_LOGIC_VECTOR(9 DOWNTO 0) := CONV_STD_LOGIC_VECTOR(92, 10);
	SIGNAL margin_y : STD_LOGIC_VECTOR(9 DOWNTO 0) := CONV_STD_LOGIC_VECTOR(4, 10);
	--MARK: signal for cells (x)
	SIGNAL cell_size : STD_LOGIC_VECTOR(9 DOWNTO 0) := CONV_STD_LOGIC_VECTOR(50, 10);
	SIGNAL cell_01x, cell_09x, cell_17x, cell_25x : STD_LOGIC_VECTOR(9 DOWNTO 0) := CONV_STD_LOGIC_VECTOR(92, 10);
	SIGNAL cell_02x, cell_10x, cell_18x, cell_26x : STD_LOGIC_VECTOR(9 DOWNTO 0) := CONV_STD_LOGIC_VECTOR(150, 10);
	SIGNAL cell_03x, cell_11x, cell_19x, cell_27x : STD_LOGIC_VECTOR(9 DOWNTO 0) := CONV_STD_LOGIC_VECTOR(208, 10);
	SIGNAL cell_04x, cell_12x, cell_20x, cell_28x : STD_LOGIC_VECTOR(9 DOWNTO 0) := CONV_STD_LOGIC_VECTOR(266, 10);
	SIGNAL cell_05x, cell_13x, cell_21x, cell_29x : STD_LOGIC_VECTOR(9 DOWNTO 0) := CONV_STD_LOGIC_VECTOR(324, 10);
	SIGNAL cell_06x, cell_14x, cell_22x, cell_30x : STD_LOGIC_VECTOR(9 DOWNTO 0) := CONV_STD_LOGIC_VECTOR(382, 10);
	SIGNAL cell_07x, cell_15x, cell_23x, cell_31x : STD_LOGIC_VECTOR(9 DOWNTO 0) := CONV_STD_LOGIC_VECTOR(440, 10);
	SIGNAL cell_08x, cell_16x, cell_24x, cell_32x : STD_LOGIC_VECTOR(9 DOWNTO 0) := CONV_STD_LOGIC_VECTOR(498, 10);
	SIGNAL cell_33x, cell_41x, cell_49x, cell_57x : STD_LOGIC_VECTOR(9 DOWNTO 0) := CONV_STD_LOGIC_VECTOR(92, 10);
	SIGNAL cell_34x, cell_42x, cell_50x, cell_58x : STD_LOGIC_VECTOR(9 DOWNTO 0) := CONV_STD_LOGIC_VECTOR(150, 10);
	SIGNAL cell_35x, cell_43x, cell_51x, cell_59x : STD_LOGIC_VECTOR(9 DOWNTO 0) := CONV_STD_LOGIC_VECTOR(208, 10);
	SIGNAL cell_36x, cell_44x, cell_52x, cell_60x : STD_LOGIC_VECTOR(9 DOWNTO 0) := CONV_STD_LOGIC_VECTOR(266, 10);
	SIGNAL cell_37x, cell_45x, cell_53x, cell_61x : STD_LOGIC_VECTOR(9 DOWNTO 0) := CONV_STD_LOGIC_VECTOR(324, 10);
	SIGNAL cell_38x, cell_46x, cell_54x, cell_62x : STD_LOGIC_VECTOR(9 DOWNTO 0) := CONV_STD_LOGIC_VECTOR(382, 10);
	SIGNAL cell_39x, cell_47x, cell_55x, cell_63x : STD_LOGIC_VECTOR(9 DOWNTO 0) := CONV_STD_LOGIC_VECTOR(440, 10);
	SIGNAL cell_40x, cell_48x, cell_56x, cell_64x : STD_LOGIC_VECTOR(9 DOWNTO 0) := CONV_STD_LOGIC_VECTOR(498, 10);
	--MARK: signal for cells (y)
	SIGNAL cell_01y, cell_02y, cell_03y, cell_04y : STD_LOGIC_VECTOR(9 DOWNTO 0) := CONV_STD_LOGIC_VECTOR(4, 10);
	SIGNAL cell_05y, cell_06y, cell_07y, cell_08y : STD_LOGIC_VECTOR(9 DOWNTO 0) := CONV_STD_LOGIC_VECTOR(4, 10);
	SIGNAL cell_09y, cell_10y, cell_11y, cell_12y : STD_LOGIC_VECTOR(9 DOWNTO 0) := CONV_STD_LOGIC_VECTOR(62, 10);
	SIGNAL cell_13y, cell_14y, cell_15y, cell_16y : STD_LOGIC_VECTOR(9 DOWNTO 0) := CONV_STD_LOGIC_VECTOR(62, 10);
	SIGNAL cell_17y, cell_18y, cell_19y, cell_20y : STD_LOGIC_VECTOR(9 DOWNTO 0) := CONV_STD_LOGIC_VECTOR(120, 10);
	SIGNAL cell_21y, cell_22y, cell_23y, cell_24y : STD_LOGIC_VECTOR(9 DOWNTO 0) := CONV_STD_LOGIC_VECTOR(120, 10);
	SIGNAL cell_25y, cell_26y, cell_27y, cell_28y : STD_LOGIC_VECTOR(9 DOWNTO 0) := CONV_STD_LOGIC_VECTOR(178, 10);
	SIGNAL cell_29y, cell_30y, cell_31y, cell_32y : STD_LOGIC_VECTOR(9 DOWNTO 0) := CONV_STD_LOGIC_VECTOR(178, 10);
	SIGNAL cell_33y, cell_34y, cell_35y, cell_36y : STD_LOGIC_VECTOR(9 DOWNTO 0) := CONV_STD_LOGIC_VECTOR(236, 10);
	SIGNAL cell_37y, cell_38y, cell_39y, cell_40y : STD_LOGIC_VECTOR(9 DOWNTO 0) := CONV_STD_LOGIC_VECTOR(236, 10);
	SIGNAL cell_41y, cell_42y, cell_43y, cell_44y : STD_LOGIC_VECTOR(9 DOWNTO 0) := CONV_STD_LOGIC_VECTOR(294, 10);
	SIGNAL cell_45y, cell_46y, cell_47y, cell_48y : STD_LOGIC_VECTOR(9 DOWNTO 0) := CONV_STD_LOGIC_VECTOR(294, 10);
	SIGNAL cell_49y, cell_50y, cell_51y, cell_52y : STD_LOGIC_VECTOR(9 DOWNTO 0) := CONV_STD_LOGIC_VECTOR(352, 10);
	SIGNAL cell_53y, cell_54y, cell_55y, cell_56y : STD_LOGIC_VECTOR(9 DOWNTO 0) := CONV_STD_LOGIC_VECTOR(352, 10);
	SIGNAL cell_57y, cell_58y, cell_59y, cell_60y : STD_LOGIC_VECTOR(9 DOWNTO 0) := CONV_STD_LOGIC_VECTOR(410, 10);
	SIGNAL cell_61y, cell_62y, cell_63y, cell_64y : STD_LOGIC_VECTOR(9 DOWNTO 0) := CONV_STD_LOGIC_VECTOR(410, 10);
	--MARK: signal for bitmaps
	TYPE number_bitmap IS ARRAY(0 TO 49, 0 TO 49) OF STD_LOGIC;
	SIGNAL number_0 : number_bitmap := (
		"00000000000000000001111111111111111110000000000000",
		"00000000000000000011111111111111111111000000000000",
		"00000000000000000111111111111111111111100000000000",
		"00000000000000011111111111111111111111110000000000",
		"00000000000000111111111111111111111111111000000000",
		"00000000000001111111111111111111111111111100000000",
		"00000000000001111111000000000000000011111100000000",
		"00000000000001111111000000000000000111111100000000",
		"00000000000001111111000000000000000111111000000000",
		"00000000000011111110000000000000000111111000000000",
		"00000000000011111110000000000000000111111000000000",
		"00000000000011111110000000000000000111111000000000",
		"00000000000011111110000000000000000111111000000000",
		"00000000000011111110000000000000001111111000000000",
		"00000000000011111110000000000000001111111000000000",
		"00000000000111111100000000000000001111110000000000",
		"00000000000111111100000000000000001111110000000000",
		"00000000000111111100000000000000001111110000000000",
		"00000000000111111100000000000000001111110000000000",
		"00000000000111111100000000000000001111110000000000",
		"00000000000111111100000000000000011111110000000000",
		"00000000000111111000000000000000011111100000000000",
		"00000000000111111111111111111111111111100000000000",
		"00000000000111110000000000000000001111000000000000",
		"00000000000011100000000000000000000110000000000000",
		"00000000000011000000000000000000000110000000000000",
		"00000000000011100000000000000000001110000000000000",
		"00000000000111111111111111111111111111000000000000",
		"00000000001111110000000000000000111111000000000000",
		"00000000001111110000000000000000111111000000000000",
		"00000000001111110000000000000000111111000000000000",
		"00000000011111110000000000000000111111000000000000",
		"00000000011111110000000000000000111111000000000000",
		"00000000011111110000000000000000111111000000000000",
		"00000000011111100000000000000001111111000000000000",
		"00000000011111100000000000000001111111000000000000",
		"00000000111111100000000000000001111110000000000000",
		"00000000111111100000000000000001111110000000000000",
		"00000000111111100000000000000001111110000000000000",
		"00000000111111100000000000000001111110000000000000",
		"00000000111111100000000000000001111110000000000000",
		"00000000111111000000000000000011111110000000000000",
		"00000000111111000000000000000011111110000000000000",
		"00000001111111000000000000000011111100000000000000",
		"00000001111111111111111111111111111100000000000000",
		"00000001111111111111111111111111111000000000000000",
		"00000000111111111111111111111111110000000000000000",
		"00000000011111111111111111111111100000000000000000",
		"00000000001111111111111111111111000000000000000000",
		"00000000000111111111111111111110000000000000000000");
	SIGNAL number_1 : number_bitmap := (
		"00000000000000000001111111111111111110000000000000",
		"00000000000000000010000000000000000001000000000000",
		"00000000000000000100000000000000000000100000000000",
		"00000000000000011100000000000000000000110000000000",
		"00000000000000100010000000000000000001111000000000",
		"00000000000001000011111111111111111111111100000000",
		"00000000000001000001000000000000000011111100000000",
		"00000000000001000001000000000000000111111100000000",
		"00000000000001000001000000000000000111111000000000",
		"00000000000010000010000000000000000111111000000000",
		"00000000000010000010000000000000000111111000000000",
		"00000000000010000010000000000000000111111000000000",
		"00000000000010000010000000000000000111111000000000",
		"00000000000010000010000000000000001111111000000000",
		"00000000000010000010000000000000001111111000000000",
		"00000000000100000100000000000000001111110000000000",
		"00000000000100000100000000000000001111110000000000",
		"00000000000100000100000000000000001111110000000000",
		"00000000000100000100000000000000001111110000000000",
		"00000000000100000100000000000000001111110000000000",
		"00000000000100000100000000000000011111110000000000",
		"00000000000100001000000000000000011111100000000000",
		"00000000000100001111111111111111111111100000000000",
		"00000000000100010000000000000000001111000000000000",
		"00000000000010100000000000000000000110000000000000",
		"00000000000011000000000000000000000110000000000000",
		"00000000000010100000000000000000001110000000000000",
		"00000000000100011111111111111111111111000000000000",
		"00000000001000010000000000000000111111000000000000",
		"00000000001000010000000000000000111111000000000000",
		"00000000001000010000000000000000111111000000000000",
		"00000000010000010000000000000000111111000000000000",
		"00000000010000010000000000000000111111000000000000",
		"00000000010000010000000000000000111111000000000000",
		"00000000010000100000000000000001111111000000000000",
		"00000000010000100000000000000001111111000000000000",
		"00000000100000100000000000000001111110000000000000",
		"00000000100000100000000000000001111110000000000000",
		"00000000100000100000000000000001111110000000000000",
		"00000000100000100000000000000001111110000000000000",
		"00000000100000100000000000000001111110000000000000",
		"00000000100001000000000000000011111110000000000000",
		"00000000100001000000000000000011111110000000000000",
		"00000001000001000000000000000011111100000000000000",
		"00000001000001111111111111111111111100000000000000",
		"00000001000010000000000000000001111000000000000000",
		"00000000100100000000000000000000110000000000000000",
		"00000000011000000000000000000000100000000000000000",
		"00000000001000000000000000000001000000000000000000",
		"00000000000111111111111111111110000000000000000000");
	SIGNAL number_2 : number_bitmap := (
		"00000000000000000001111111111111111110000000000000",
		"00000000000000000011111111111111111111000000000000",
		"00000000000000000111111111111111111111100000000000",
		"00000000000000011111111111111111111111110000000000",
		"00000000000000100011111111111111111111111000000000",
		"00000000000001000011111111111111111111111100000000",
		"00000000000001000001000000000000000011111100000000",
		"00000000000001000001000000000000000111111100000000",
		"00000000000001000001000000000000000111111000000000",
		"00000000000010000010000000000000000111111000000000",
		"00000000000010000010000000000000000111111000000000",
		"00000000000010000010000000000000000111111000000000",
		"00000000000010000010000000000000000111111000000000",
		"00000000000010000010000000000000001111111000000000",
		"00000000000010000010000000000000001111111000000000",
		"00000000000100000100000000000000001111110000000000",
		"00000000000100000100000000000000001111110000000000",
		"00000000000100000100000000000000001111110000000000",
		"00000000000100000100000000000000001111110000000000",
		"00000000000100000100000000000000001111110000000000",
		"00000000000100000100000000000000011111110000000000",
		"00000000000100001000000000000000011111100000000000",
		"00000000000100001111111111111111111111100000000000",
		"00000000000100011111111111111111111111000000000000",
		"00000000000010111111111111111111111110000000000000",
		"00000000000011111111111111111111111110000000000000",
		"00000000000011111111111111111111111010000000000000",
		"00000000000111111111111111111111110001000000000000",
		"00000000001111110000000000000000100001000000000000",
		"00000000001111110000000000000000100001000000000000",
		"00000000001111110000000000000000100001000000000000",
		"00000000011111110000000000000000100001000000000000",
		"00000000011111110000000000000000100001000000000000",
		"00000000011111110000000000000000100001000000000000",
		"00000000011111100000000000000001000001000000000000",
		"00000000011111100000000000000001000001000000000000",
		"00000000111111100000000000000001000010000000000000",
		"00000000111111100000000000000001000010000000000000",
		"00000000111111100000000000000001000010000000000000",
		"00000000111111100000000000000001000010000000000000",
		"00000000111111100000000000000001000010000000000000",
		"00000000111111000000000000000010000010000000000000",
		"00000000111111000000000000000010000010000000000000",
		"00000001111111000000000000000010000100000000000000",
		"00000001111111111111111111111110000100000000000000",
		"00000001111111111111111111111111001000000000000000",
		"00000000111111111111111111111111110000000000000000",
		"00000000011111111111111111111111100000000000000000",
		"00000000001111111111111111111111000000000000000000",
		"00000000000111111111111111111110000000000000000000");
	SIGNAL number_3 : number_bitmap := (
		"00000000000000000001111111111111111110000000000000",
		"00000000000000000011111111111111111111000000000000",
		"00000000000000000111111111111111111111100000000000",
		"00000000000000011111111111111111111111110000000000",
		"00000000000000100011111111111111111111111000000000",
		"00000000000001000011111111111111111111111100000000",
		"00000000000001000001000000000000000011111100000000",
		"00000000000001000001000000000000000111111100000000",
		"00000000000001000001000000000000000111111000000000",
		"00000000000010000010000000000000000111111000000000",
		"00000000000010000010000000000000000111111000000000",
		"00000000000010000010000000000000000111111000000000",
		"00000000000010000010000000000000000111111000000000",
		"00000000000010000010000000000000001111111000000000",
		"00000000000010000010000000000000001111111000000000",
		"00000000000100000100000000000000001111110000000000",
		"00000000000100000100000000000000001111110000000000",
		"00000000000100000100000000000000001111110000000000",
		"00000000000100000100000000000000001111110000000000",
		"00000000000100000100000000000000001111110000000000",
		"00000000000100000100000000000000011111110000000000",
		"00000000000100001000000000000000011111100000000000",
		"00000000000100001111111111111111111111100000000000",
		"00000000000100011111111111111111111111000000000000",
		"00000000000010111111111111111111111110000000000000",
		"00000000000011111111111111111111111110000000000000",
		"00000000000010111111111111111111111110000000000000",
		"00000000000100011111111111111111111111000000000000",
		"00000000001000010000000000000000111111000000000000",
		"00000000001000010000000000000000111111000000000000",
		"00000000001000010000000000000000111111000000000000",
		"00000000010000010000000000000000111111000000000000",
		"00000000010000010000000000000000111111000000000000",
		"00000000010000010000000000000000111111000000000000",
		"00000000010000100000000000000001111111000000000000",
		"00000000010000100000000000000001111111000000000000",
		"00000000100000100000000000000001111110000000000000",
		"00000000100000100000000000000001111110000000000000",
		"00000000100000100000000000000001111110000000000000",
		"00000000100000100000000000000001111110000000000000",
		"00000000100000100000000000000001111110000000000000",
		"00000000100001000000000000000011111110000000000000",
		"00000000100001000000000000000011111110000000000000",
		"00000001000001000000000000000011111100000000000000",
		"00000001000001111111111111111111111100000000000000",
		"00000001000011111111111111111111111000000000000000",
		"00000000100111111111111111111111110000000000000000",
		"00000000011111111111111111111111100000000000000000",
		"00000000001111111111111111111111000000000000000000",
		"00000000000111111111111111111110000000000000000000");
	SIGNAL number_4 : number_bitmap := (
		"00000000000000000001111111111111111110000000000000",
		"00000000000000000010000000000000000001000000000000",
		"00000000000000000100000000000000000000100000000000",
		"00000000000000011100000000000000000000110000000000",
		"00000000000000111110000000000000000001111000000000",
		"00000000000001111111111111111111111111111100000000",
		"00000000000001111111000000000000000011111100000000",
		"00000000000001111111000000000000000111111100000000",
		"00000000000001111111000000000000000111111000000000",
		"00000000000011111110000000000000000111111000000000",
		"00000000000011111110000000000000000111111000000000",
		"00000000000011111110000000000000000111111000000000",
		"00000000000011111110000000000000000111111000000000",
		"00000000000011111110000000000000001111111000000000",
		"00000000000011111110000000000000001111111000000000",
		"00000000000111111100000000000000001111110000000000",
		"00000000000111111100000000000000001111110000000000",
		"00000000000111111100000000000000001111110000000000",
		"00000000000111111100000000000000001111110000000000",
		"00000000000111111100000000000000001111110000000000",
		"00000000000111111100000000000000011111110000000000",
		"00000000000111111000000000000000011111100000000000",
		"00000000000111111111111111111111111111100000000000",
		"00000000000111111111111111111111111111000000000000",
		"00000000000011111111111111111111111110000000000000",
		"00000000000011111111111111111111111110000000000000",
		"00000000000010111111111111111111111110000000000000",
		"00000000000100011111111111111111111111000000000000",
		"00000000001000010000000000000000111111000000000000",
		"00000000001000010000000000000000111111000000000000",
		"00000000001000010000000000000000111111000000000000",
		"00000000010000010000000000000000111111000000000000",
		"00000000010000010000000000000000111111000000000000",
		"00000000010000010000000000000000111111000000000000",
		"00000000010000100000000000000001111111000000000000",
		"00000000010000100000000000000001111111000000000000",
		"00000000100000100000000000000001111110000000000000",
		"00000000100000100000000000000001111110000000000000",
		"00000000100000100000000000000001111110000000000000",
		"00000000100000100000000000000001111110000000000000",
		"00000000100000100000000000000001111110000000000000",
		"00000000100001000000000000000011111110000000000000",
		"00000000100001000000000000000011111110000000000000",
		"00000001000001000000000000000011111100000000000000",
		"00000001000001111111111111111111111100000000000000",
		"00000001000010000000000000000001111000000000000000",
		"00000000100100000000000000000000110000000000000000",
		"00000000011000000000000000000000100000000000000000",
		"00000000001000000000000000000001000000000000000000",
		"00000000000111111111111111111110000000000000000000");
	SIGNAL number_5 : number_bitmap := (
		"00000000000000000001111111111111111110000000000000",
		"00000000000000000011111111111111111111000000000000",
		"00000000000000000111111111111111111111100000000000",
		"00000000000000011111111111111111111111110000000000",
		"00000000000000111111111111111111111111001000000000",
		"00000000000001111111111111111111111110000100000000",
		"00000000000001111111000000000000000010000100000000",
		"00000000000001111111000000000000000100001100000000",
		"00000000000001111111000000000000000100001000000000",
		"00000000000011111110000000000000000100001000000000",
		"00000000000011111110000000000000000100001000000000",
		"00000000000011111110000000000000000100001000000000",
		"00000000000011111110000000000000000100001000000000",
		"00000000000011111110000000000000001000001000000000",
		"00000000000011111110000000000000001000001000000000",
		"00000000000111111100000000000000001000010000000000",
		"00000000000111111100000000000000001000010000000000",
		"00000000000111111100000000000000001000010000000000",
		"00000000000111111100000000000000001000010000000000",
		"00000000000111111100000000000000001000010000000000",
		"00000000000111111100000000000000010000010000000000",
		"00000000000111111000000000000000010000100000000000",
		"00000000000111111111111111111111110000100000000000",
		"00000000000111111111111111111111111001000000000000",
		"00000000000011111111111111111111111110000000000000",
		"00000000000011111111111111111111111110000000000000",
		"00000000000010111111111111111111111110000000000000",
		"00000000000100011111111111111111111111000000000000",
		"00000000001000010000000000000000111111000000000000",
		"00000000001000010000000000000000111111000000000000",
		"00000000001000010000000000000000111111000000000000",
		"00000000010000010000000000000000111111000000000000",
		"00000000010000010000000000000000111111000000000000",
		"00000000010000010000000000000000111111000000000000",
		"00000000010000100000000000000001111111000000000000",
		"00000000010000100000000000000001111111000000000000",
		"00000000100000100000000000000001111110000000000000",
		"00000000100000100000000000000001111110000000000000",
		"00000000100000100000000000000001111110000000000000",
		"00000000100000100000000000000001111110000000000000",
		"00000000100000100000000000000001111110000000000000",
		"00000000100001000000000000000011111110000000000000",
		"00000000100001000000000000000011111110000000000000",
		"00000001000001000000000000000011111100000000000000",
		"00000001000001111111111111111111111100000000000000",
		"00000001000011111111111111111111111000000000000000",
		"00000000100111111111111111111111110000000000000000",
		"00000000011111111111111111111111100000000000000000",
		"00000000001111111111111111111111000000000000000000",
		"00000000000111111111111111111110000000000000000000");
	SIGNAL number_6 : number_bitmap := (
		"00000000000000000001111111111111111110000000000000",
		"00000000000000000011111111111111111111000000000000",
		"00000000000000000111111111111111111111100000000000",
		"00000000000000011111111111111111111111110000000000",
		"00000000000000111111111111111111111111001000000000",
		"00000000000001111111111111111111111110000100000000",
		"00000000000001111111000000000000000010000100000000",
		"00000000000001111111000000000000000100001100000000",
		"00000000000001111111000000000000000100001000000000",
		"00000000000011111110000000000000000100001000000000",
		"00000000000011111110000000000000000100001000000000",
		"00000000000011111110000000000000000100001000000000",
		"00000000000011111110000000000000000100001000000000",
		"00000000000011111110000000000000001000001000000000",
		"00000000000011111110000000000000001000001000000000",
		"00000000000111111100000000000000001000010000000000",
		"00000000000111111100000000000000001000010000000000",
		"00000000000111111100000000000000001000010000000000",
		"00000000000111111100000000000000001000010000000000",
		"00000000000111111100000000000000001000010000000000",
		"00000000000111111100000000000000010000010000000000",
		"00000000000111111000000000000000010000100000000000",
		"00000000000111111111111111111111110000100000000000",
		"00000000000111111111111111111111111001000000000000",
		"00000000000011111111111111111111111110000000000000",
		"00000000000011111111111111111111111110000000000000",
		"00000000000011111111111111111111111110000000000000",
		"00000000000111111111111111111111111111000000000000",
		"00000000001111110000000000000000111111000000000000",
		"00000000001111110000000000000000111111000000000000",
		"00000000001111110000000000000000111111000000000000",
		"00000000011111110000000000000000111111000000000000",
		"00000000011111110000000000000000111111000000000000",
		"00000000011111110000000000000000111111000000000000",
		"00000000011111100000000000000001111111000000000000",
		"00000000011111100000000000000001111111000000000000",
		"00000000111111100000000000000001111110000000000000",
		"00000000111111100000000000000001111110000000000000",
		"00000000111111100000000000000001111110000000000000",
		"00000000111111100000000000000001111110000000000000",
		"00000000111111100000000000000001111110000000000000",
		"00000000111111000000000000000011111110000000000000",
		"00000000111111000000000000000011111110000000000000",
		"00000001111111000000000000000011111100000000000000",
		"00000001111111111111111111111111111100000000000000",
		"00000001111111111111111111111111111000000000000000",
		"00000000111111111111111111111111110000000000000000",
		"00000000011111111111111111111111100000000000000000",
		"00000000001111111111111111111111000000000000000000",
		"00000000000111111111111111111110000000000000000000");
	SIGNAL number_7 : number_bitmap := (
		"00000000000000000001111111111111111110000000000000",
		"00000000000000000011111111111111111111000000000000",
		"00000000000000000111111111111111111111100000000000",
		"00000000000000011111111111111111111111110000000000",
		"00000000000000100011111111111111111111111000000000",
		"00000000000001000011111111111111111111111100000000",
		"00000000000001000001000000000000000011111100000000",
		"00000000000001000001000000000000000111111100000000",
		"00000000000001000001000000000000000111111000000000",
		"00000000000010000010000000000000000111111000000000",
		"00000000000010000010000000000000000111111000000000",
		"00000000000010000010000000000000000111111000000000",
		"00000000000010000010000000000000000111111000000000",
		"00000000000010000010000000000000001111111000000000",
		"00000000000010000010000000000000001111111000000000",
		"00000000000100000100000000000000001111110000000000",
		"00000000000100000100000000000000001111110000000000",
		"00000000000100000100000000000000001111110000000000",
		"00000000000100000100000000000000001111110000000000",
		"00000000000100000100000000000000001111110000000000",
		"00000000000100000100000000000000011111110000000000",
		"00000000000100001000000000000000011111100000000000",
		"00000000000100001111111111111111111111100000000000",
		"00000000000100010000000000000000001111000000000000",
		"00000000000010100000000000000000000110000000000000",
		"00000000000011000000000000000000000110000000000000",
		"00000000000010100000000000000000001110000000000000",
		"00000000000100011111111111111111111111000000000000",
		"00000000001000010000000000000000111111000000000000",
		"00000000001000010000000000000000111111000000000000",
		"00000000001000010000000000000000111111000000000000",
		"00000000010000010000000000000000111111000000000000",
		"00000000010000010000000000000000111111000000000000",
		"00000000010000010000000000000000111111000000000000",
		"00000000010000100000000000000001111111000000000000",
		"00000000010000100000000000000001111111000000000000",
		"00000000100000100000000000000001111110000000000000",
		"00000000100000100000000000000001111110000000000000",
		"00000000100000100000000000000001111110000000000000",
		"00000000100000100000000000000001111110000000000000",
		"00000000100000100000000000000001111110000000000000",
		"00000000100001000000000000000011111110000000000000",
		"00000000100001000000000000000011111110000000000000",
		"00000001000001000000000000000011111100000000000000",
		"00000001000001111111111111111111111100000000000000",
		"00000001000010000000000000000001111000000000000000",
		"00000000100100000000000000000000110000000000000000",
		"00000000011000000000000000000000100000000000000000",
		"00000000001000000000000000000001000000000000000000",
		"00000000000111111111111111111110000000000000000000");
	SIGNAL number_8 : number_bitmap := (
		"00000000000000000001111111111111111110000000000000",
		"00000000000000000011111111111111111111000000000000",
		"00000000000000000111111111111111111111100000000000",
		"00000000000000011111111111111111111111110000000000",
		"00000000000000111111111111111111111111111000000000",
		"00000000000001111111111111111111111111111100000000",
		"00000000000001111111000000000000000011111100000000",
		"00000000000001111111000000000000000111111100000000",
		"00000000000001111111000000000000000111111000000000",
		"00000000000011111110000000000000000111111000000000",
		"00000000000011111110000000000000000111111000000000",
		"00000000000011111110000000000000000111111000000000",
		"00000000000011111110000000000000000111111000000000",
		"00000000000011111110000000000000001111111000000000",
		"00000000000011111110000000000000001111111000000000",
		"00000000000111111100000000000000001111110000000000",
		"00000000000111111100000000000000001111110000000000",
		"00000000000111111100000000000000001111110000000000",
		"00000000000111111100000000000000001111110000000000",
		"00000000000111111100000000000000001111110000000000",
		"00000000000111111100000000000000011111110000000000",
		"00000000000111111000000000000000011111100000000000",
		"00000000000111111111111111111111111111100000000000",
		"00000000000111111111111111111111111111000000000000",
		"00000000000011111111111111111111111110000000000000",
		"00000000000011111111111111111111111110000000000000",
		"00000000000011111111111111111111111110000000000000",
		"00000000000111111111111111111111111111000000000000",
		"00000000001111110000000000000000111111000000000000",
		"00000000001111110000000000000000111111000000000000",
		"00000000001111110000000000000000111111000000000000",
		"00000000011111110000000000000000111111000000000000",
		"00000000011111110000000000000000111111000000000000",
		"00000000011111110000000000000000111111000000000000",
		"00000000011111100000000000000001111111000000000000",
		"00000000011111100000000000000001111111000000000000",
		"00000000111111100000000000000001111110000000000000",
		"00000000111111100000000000000001111110000000000000",
		"00000000111111100000000000000001111110000000000000",
		"00000000111111100000000000000001111110000000000000",
		"00000000111111100000000000000001111110000000000000",
		"00000000111111000000000000000011111110000000000000",
		"00000000111111000000000000000011111110000000000000",
		"00000001111111000000000000000011111100000000000000",
		"00000001111111111111111111111111111100000000000000",
		"00000001111111111111111111111111111000000000000000",
		"00000000111111111111111111111111110000000000000000",
		"00000000011111111111111111111111100000000000000000",
		"00000000001111111111111111111111000000000000000000",
		"00000000000111111111111111111110000000000000000000");
	SIGNAL number_empty : number_bitmap := (
		"00000000000000000001111111111111111110000000000000",
		"00000000000000000010000000000000000001000000000000",
		"00000000000000000100000000000000000000100000000000",
		"00000000000000011100000000000000000000110000000000",
		"00000000000000100010000000000000000001001000000000",
		"00000000000001000011111111111111111110000100000000",
		"00000000000001000001000000000000000010000100000000",
		"00000000000001000001000000000000000100001100000000",
		"00000000000001000001000000000000000100001000000000",
		"00000000000010000010000000000000000100001000000000",
		"00000000000010000010000000000000000100001000000000",
		"00000000000010000010000000000000000100001000000000",
		"00000000000010000010000000000000000100001000000000",
		"00000000000010000010000000000000001000001000000000",
		"00000000000010000010000000000000001000001000000000",
		"00000000000100000100000000000000001000010000000000",
		"00000000000100000100000000000000001000010000000000",
		"00000000000100000100000000000000001000010000000000",
		"00000000000100000100000000000000001000010000000000",
		"00000000000100000100000000000000001000010000000000",
		"00000000000100000100000000000000010000010000000000",
		"00000000000100001000000000000000010000100000000000",
		"00000000000100001111111111111111110000100000000000",
		"00000000000100010000000000000000001001000000000000",
		"00000000000010100000000000000000000110000000000000",
		"00000000000011000000000000000000000110000000000000",
		"00000000000010100000000000000000001010000000000000",
		"00000000000100011111111111111111110001000000000000",
		"00000000001000010000000000000000100001000000000000",
		"00000000001000010000000000000000100001000000000000",
		"00000000001000010000000000000000100001000000000000",
		"00000000010000010000000000000000100001000000000000",
		"00000000010000010000000000000000100001000000000000",
		"00000000010000010000000000000000100001000000000000",
		"00000000010000100000000000000001000001000000000000",
		"00000000010000100000000000000001000001000000000000",
		"00000000100000100000000000000001000010000000000000",
		"00000000100000100000000000000001000010000000000000",
		"00000000100000100000000000000001000010000000000000",
		"00000000100000100000000000000001000010000000000000",
		"00000000100000100000000000000001000010000000000000",
		"00000000100001000000000000000010000010000000000000",
		"00000000100001000000000000000010000010000000000000",
		"00000001000001000000000000000010000100000000000000",
		"00000001000001111111111111111110000100000000000000",
		"00000001000010000000000000000001001000000000000000",
		"00000000100100000000000000000000110000000000000000",
		"00000000011000000000000000000000100000000000000000",
		"00000000001000000000000000000001000000000000000000",
		"00000000000111111111111111111110000000000000000000");

	PROCEDURE CellDisplay (
		cell_x : IN INTEGER;
		cell_y : IN INTEGER
	) IS
		VARIABLE pos_y : INTEGER;
		VARIABLE pos_x : INTEGER;
	BEGIN
		IF cell_status(cell_x, cell_y) = 0 THEN -- closed cell
			IF cell_flagged(cell_x, cell_y) = 0 THEN -- not flagged (green) 
				Red <= closed_cell_color(2);
				Green <= closed_cell_color(1);
				Blue <= closed_cell_color(0);
			ELSE -- flagged (red)
				Red <= flagged_cell_color(2);
				Green <= flagged_cell_color(1);
				Blue <= flagged_cell_color(0);
			END IF;
		ELSE -- open cell (black)
			pos_x := CONV_INTEGER(pixel_column - cell_08x);
			pos_y := CONV_INTEGER(pixel_row - cell_08y);

			CASE cell_value(cell_x, cell_y) IS
				WHEN 0 =>
					IF number_0(pos_y, pos_x) = '1' THEN
						Red <= opened_cell_color(2);
						Green <= opened_cell_color(1);
						Blue <= opened_cell_color(0);
					ELSE
						Red <= background_color(2);
						Green <= background_color(1);
						Blue <= background_color(0);
					END IF;
				WHEN 1 =>
					IF number_1(pos_y, pos_x) = '1' THEN
						Red <= opened_cell_color(2);
						Green <= opened_cell_color(1);
						Blue <= opened_cell_color(0);
					ELSE
						Red <= background_color(2);
						Green <= background_color(1);
						Blue <= background_color(0);
					END IF;
				WHEN 2 =>
					IF number_2(pos_y, pos_x) = '1' THEN
						Red <= opened_cell_color(2);
						Green <= opened_cell_color(1);
						Blue <= opened_cell_color(0);
					ELSE
						Red <= background_color(2);
						Green <= background_color(1);
						Blue <= background_color(0);
					END IF;
				WHEN 3 =>
					IF number_3(pos_y, pos_x) = '1' THEN
						Red <= opened_cell_color(2);
						Green <= opened_cell_color(1);
						Blue <= opened_cell_color(0);
					ELSE
						Red <= background_color(2);
						Green <= background_color(1);
						Blue <= background_color(0);
					END IF;
				WHEN 4 =>
					IF number_4(pos_y, pos_x) = '1' THEN
						Red <= opened_cell_color(2);
						Green <= opened_cell_color(1);
						Blue <= opened_cell_color(0);
					ELSE
						Red <= background_color(2);
						Green <= background_color(1);
						Blue <= background_color(0);
					END IF;
				WHEN 5 =>
					IF number_5(pos_y, pos_x) = '1' THEN
						Red <= opened_cell_color(2);
						Green <= opened_cell_color(1);
						Blue <= opened_cell_color(0);
					ELSE
						Red <= background_color(2);
						Green <= background_color(1);
						Blue <= background_color(0);
					END IF;
				WHEN 6 =>
					IF number_6(pos_y, pos_x) = '1' THEN
						Red <= opened_cell_color(2);
						Green <= opened_cell_color(1);
						Blue <= opened_cell_color(0);
					ELSE
						Red <= background_color(2);
						Green <= background_color(1);
						Blue <= background_color(0);
					END IF;
				WHEN 7 =>
					IF number_7(pos_y, pos_x) = '1' THEN
						Red <= opened_cell_color(2);
						Green <= opened_cell_color(1);
						Blue <= opened_cell_color(0);
					ELSE
						Red <= background_color(2);
						Green <= background_color(1);
						Blue <= background_color(0);
					END IF;
				WHEN 8 =>
					IF number_8(pos_y, pos_x) = '1' THEN
						Red <= opened_cell_color(2);
						Green <= opened_cell_color(1);
						Blue <= opened_cell_color(0);
					ELSE
						Red <= background_color(2);
						Green <= background_color(1);
						Blue <= background_color(0);
					END IF;
				WHEN OTHERS =>
					IF number_empty(pos_y, pos_x) = '1' THEN
						Red <= opened_cell_color(2);
						Green <= opened_cell_color(1);
						Blue <= opened_cell_color(0);
					ELSE
						Red <= background_color(2);
						Green <= background_color(1);
						Blue <= background_color(0);
					END IF;
			END CASE;
		END IF;
		-- Teyon made user position show as magenta (overrides showing flag like this)
		IF cell_x = cell_userb(0) and cell_y = cell_userb(1) then
			Red <= '1';
			Green <= '0';
			Blue <= '1';
		end if;
	END CellDisplay;
BEGIN
	--MARK: Process
	-- display the grid of the board
	RGB_Display : PROCESS (pixel_row, pixel_column)
		-- calculate the position within the bitmap

	BEGIN
		-- if-else statement (first long section is not needed <- square, not circle)
		IF -- set the background
			-- TODO: check this background color logic
			-- 1.
			(pixel_column < margin_x) AND
			(pixel_column > margin_x + margin_width) AND
			(pixel_row < margin_y) AND
			(pixel_row > margin_y + margin_height)
			-- -- 2.
			-- ('0' & pixel_column < 92) AND ('0' & pixel_column > 548) AND
			-- ('0' & pixel_row < 4) AND ('0' & pixel_row > 475)
			-- -- 3.
			-- ('0' & pixel_column < cell_01x) AND ('0' & pixel_column >= display_width - cell_01x) AND
			-- ('0' & pixel_row < cell_01y) AND ('0' & pixel_row > display_height - cell_01y)
			THEN
			-- 'background color' to white
			Red <= background_color(2);
			Green <= background_color(1);
			Blue <= background_color(0);
		ELSE -- if chains <- cell region
			IF --TODO: check this w/ & w/o `'0' &``
				-- 1.
				(cell_01x <= pixel_column) AND (pixel_column < cell_01x + cell_size) AND
				(cell_01y <= pixel_row) AND (pixel_row < cell_01y + cell_size)
				-- -- 2.
				-- ('0' & cell_01x <= pixel_column) AND ('0' & pixel_column < cell_01x + cell_size) AND
				-- ('0' & cell_01y <= pixel_row) AND ('0' & pixel_row < cell_01y + cell_size)
				-- -- 3.
				-- ('0' & pixel_column >= cell_01x) AND ('0' & pixel_column < cell_01x + cell_size) AND
				-- ('0' & pixel_row >= cell_01y) AND ('0' & pixel_row < cell_01y + cell_size)
				THEN
				CellDisplay(0, 0);
			ELSIF
				('0' & cell_02x <= pixel_column) AND ('0' & pixel_column <= cell_02x + cell_size) AND
				('0' & cell_02y <= pixel_row) AND ('0' & pixel_row <= cell_02y + cell_size)
				THEN
				CellDisplay(0, 1);
			ELSIF
				('0' & cell_03x <= pixel_column) AND ('0' & pixel_column <= cell_03x + cell_size) AND
				('0' & cell_03y <= pixel_row) AND ('0' & pixel_row <= cell_03y + cell_size)
				THEN
				CellDisplay(0, 2);
			ELSIF
				('0' & cell_04x <= pixel_column) AND ('0' & pixel_column <= cell_04x + cell_size) AND
				('0' & cell_04y <= pixel_row) AND ('0' & pixel_row <= cell_04y + cell_size)
				THEN
				CellDisplay(0, 3);
			ELSIF
				('0' & cell_05x <= pixel_column) AND ('0' & pixel_column <= cell_05x + cell_size) AND
				('0' & cell_05y <= pixel_row) AND ('0' & pixel_row <= cell_05y + cell_size)
				THEN
				CellDisplay(0, 4);
			ELSIF
				('0' & cell_06x <= pixel_column) AND ('0' & pixel_column <= cell_06x + cell_size) AND
				('0' & cell_06y <= pixel_row) AND ('0' & pixel_row <= cell_06y + cell_size)
				THEN
				CellDisplay(0, 5);
			ELSIF
				('0' & cell_07x <= pixel_column) AND ('0' & pixel_column <= cell_07x + cell_size) AND
				('0' & cell_07y <= pixel_row) AND ('0' & pixel_row <= cell_07y + cell_size)
				THEN
				CellDisplay(0, 6);
			ELSIF
				('0' & cell_08x <= pixel_column) AND ('0' & pixel_column <= cell_08x + cell_size) AND
				('0' & cell_08y <= pixel_row) AND ('0' & pixel_row <= cell_08y + cell_size)
				THEN
				CellDisplay(0, 7);
			ELSIF
				('0' & cell_09x <= pixel_column) AND ('0' & pixel_column <= cell_09x + cell_size) AND
				('0' & cell_09y <= pixel_row) AND ('0' & pixel_row <= cell_09y + cell_size)
				THEN
				CellDisplay(1, 0);
			ELSIF
				('0' & cell_10x <= pixel_column) AND ('0' & pixel_column <= cell_10x + cell_size) AND
				('0' & cell_10y <= pixel_row) AND ('0' & pixel_row <= cell_10y + cell_size)
				THEN
				CellDisplay(1, 1);
			ELSIF
				('0' & cell_11x <= pixel_column) AND ('0' & pixel_column <= cell_11x + cell_size) AND
				('0' & cell_11y <= pixel_row) AND ('0' & pixel_row <= cell_11y + cell_size)
				THEN
				CellDisplay(1, 2);
			ELSIF
				('0' & cell_12x <= pixel_column) AND ('0' & pixel_column <= cell_12x + cell_size) AND
				('0' & cell_12y <= pixel_row) AND ('0' & pixel_row <= cell_12y + cell_size)
				THEN
				CellDisplay(1, 3);
			ELSIF
				('0' & cell_13x <= pixel_column) AND ('0' & pixel_column <= cell_13x + cell_size) AND
				('0' & cell_13y <= pixel_row) AND ('0' & pixel_row <= cell_13y + cell_size)
				THEN
				CellDisplay(1, 4);
			ELSIF
				('0' & cell_14x <= pixel_column) AND ('0' & pixel_column <= cell_14x + cell_size) AND
				('0' & cell_14y <= pixel_row) AND ('0' & pixel_row <= cell_14y + cell_size)
				THEN
				CellDisplay(1, 5);
			ELSIF
				('0' & cell_15x <= pixel_column) AND ('0' & pixel_column <= cell_15x + cell_size) AND
				('0' & cell_15y <= pixel_row) AND ('0' & pixel_row <= cell_15y + cell_size)
				THEN
				CellDisplay(1, 6);
			ELSIF
				('0' & cell_16x <= pixel_column) AND ('0' & pixel_column <= cell_16x + cell_size) AND
				('0' & cell_16y <= pixel_row) AND ('0' & pixel_row <= cell_16y + cell_size)
				THEN
				CellDisplay(1, 7);
			ELSIF
				('0' & cell_17x <= pixel_column) AND ('0' & pixel_column <= cell_17x + cell_size) AND
				('0' & cell_17y <= pixel_row) AND ('0' & pixel_row <= cell_17y + cell_size)
				THEN
				CellDisplay(2, 0);
			ELSIF
				('0' & cell_18x <= pixel_column) AND ('0' & pixel_column <= cell_18x + cell_size) AND
				('0' & cell_18y <= pixel_row) AND ('0' & pixel_row <= cell_18y + cell_size)
				THEN
				CellDisplay(2, 1);
			ELSIF
				('0' & cell_19x <= pixel_column) AND ('0' & pixel_column <= cell_19x + cell_size) AND
				('0' & cell_19y <= pixel_row) AND ('0' & pixel_row <= cell_19y + cell_size)
				THEN
				CellDisplay(2, 2);
			ELSIF
				('0' & cell_20x <= pixel_column) AND ('0' & pixel_column <= cell_20x + cell_size) AND
				('0' & cell_20y <= pixel_row) AND ('0' & pixel_row <= cell_20y + cell_size)
				THEN
				CellDisplay(2, 3);
			ELSIF
				('0' & cell_21x <= pixel_column) AND ('0' & pixel_column <= cell_21x + cell_size) AND
				('0' & cell_21y <= pixel_row) AND ('0' & pixel_row <= cell_21y + cell_size)
				THEN
				CellDisplay(2, 4);
			ELSIF
				('0' & cell_22x <= pixel_column) AND ('0' & pixel_column <= cell_22x + cell_size) AND
				('0' & cell_22y <= pixel_row) AND ('0' & pixel_row <= cell_22y + cell_size)
				THEN
				CellDisplay(2, 5);
			ELSIF
				('0' & cell_23x <= pixel_column) AND ('0' & pixel_column <= cell_23x + cell_size) AND
				('0' & cell_23y <= pixel_row) AND ('0' & pixel_row <= cell_23y + cell_size)
				THEN
				CellDisplay(2, 6);
			ELSIF
				('0' & cell_24x <= pixel_column) AND ('0' & pixel_column <= cell_24x + cell_size) AND
				('0' & cell_24y <= pixel_row) AND ('0' & pixel_row <= cell_24y + cell_size)
				THEN
				CellDisplay(2, 7);
			ELSIF
				('0' & cell_25x <= pixel_column) AND ('0' & pixel_column <= cell_25x + cell_size) AND
				('0' & cell_25y <= pixel_row) AND ('0' & pixel_row <= cell_25y + cell_size)
				THEN
				CellDisplay(3, 0);
			ELSIF
				('0' & cell_26x <= pixel_column) AND ('0' & pixel_column <= cell_26x + cell_size) AND
				('0' & cell_26y <= pixel_row) AND ('0' & pixel_row <= cell_26y + cell_size)
				THEN
				CellDisplay(3, 1);
			ELSIF
				('0' & cell_27x <= pixel_column) AND ('0' & pixel_column <= cell_27x + cell_size) AND
				('0' & cell_27y <= pixel_row) AND ('0' & pixel_row <= cell_27y + cell_size)
				THEN
				CellDisplay(3, 2);
			ELSIF
				('0' & cell_28x <= pixel_column) AND ('0' & pixel_column <= cell_28x + cell_size) AND
				('0' & cell_28y <= pixel_row) AND ('0' & pixel_row <= cell_28y + cell_size)
				THEN
				CellDisplay(3, 3);
			ELSIF
				('0' & cell_29x <= pixel_column) AND ('0' & pixel_column <= cell_29x + cell_size) AND
				('0' & cell_29y <= pixel_row) AND ('0' & pixel_row <= cell_29y + cell_size)
				THEN
				CellDisplay(3, 4);
			ELSIF
				('0' & cell_30x <= pixel_column) AND ('0' & pixel_column <= cell_30x + cell_size) AND
				('0' & cell_30y <= pixel_row) AND ('0' & pixel_row <= cell_30y + cell_size)
				THEN
				CellDisplay(3, 5);
			ELSIF
				('0' & cell_31x <= pixel_column) AND ('0' & pixel_column <= cell_31x + cell_size) AND
				('0' & cell_31y <= pixel_row) AND ('0' & pixel_row <= cell_31y + cell_size)
				THEN
				CellDisplay(3, 6);
			ELSIF
				('0' & cell_32x <= pixel_column) AND ('0' & pixel_column <= cell_32x + cell_size) AND
				('0' & cell_32y <= pixel_row) AND ('0' & pixel_row <= cell_32y + cell_size)
				THEN
				CellDisplay(3, 7);
			ELSIF
				('0' & cell_33x <= pixel_column) AND ('0' & pixel_column <= cell_33x + cell_size) AND
				('0' & cell_33y <= pixel_row) AND ('0' & pixel_row <= cell_33y + cell_size)
				THEN
				CellDisplay(4, 0);
			ELSIF
				('0' & cell_34x <= pixel_column) AND ('0' & pixel_column <= cell_34x + cell_size) AND
				('0' & cell_34y <= pixel_row) AND ('0' & pixel_row <= cell_34y + cell_size)
				THEN
				CellDisplay(4, 1);
			ELSIF
				('0' & cell_35x <= pixel_column) AND ('0' & pixel_column <= cell_35x + cell_size) AND
				('0' & cell_35y <= pixel_row) AND ('0' & pixel_row <= cell_35y + cell_size)
				THEN
				CellDisplay(4, 2);
			ELSIF
				('0' & cell_36x <= pixel_column) AND ('0' & pixel_column <= cell_36x + cell_size) AND
				('0' & cell_36y <= pixel_row) AND ('0' & pixel_row <= cell_36y + cell_size)
				THEN
				CellDisplay(4, 3);
			ELSIF
				('0' & cell_37x <= pixel_column) AND ('0' & pixel_column <= cell_37x + cell_size) AND
				('0' & cell_37y <= pixel_row) AND ('0' & pixel_row <= cell_37y + cell_size)
				THEN
				CellDisplay(4, 4);
			ELSIF
				('0' & cell_38x <= pixel_column) AND ('0' & pixel_column <= cell_38x + cell_size) AND
				('0' & cell_38y <= pixel_row) AND ('0' & pixel_row <= cell_38y + cell_size)
				THEN
				CellDisplay(4, 5);
			ELSIF
				('0' & cell_39x <= pixel_column) AND ('0' & pixel_column <= cell_39x + cell_size) AND
				('0' & cell_39y <= pixel_row) AND ('0' & pixel_row <= cell_39y + cell_size)
				THEN
				CellDisplay(4, 6);
			ELSIF
				('0' & cell_40x <= pixel_column) AND ('0' & pixel_column <= cell_40x + cell_size) AND
				('0' & cell_40y <= pixel_row) AND ('0' & pixel_row <= cell_40y + cell_size)
				THEN
				CellDisplay(4, 7);
			ELSIF
				('0' & cell_41x <= pixel_column) AND ('0' & pixel_column <= cell_41x + cell_size) AND
				('0' & cell_41y <= pixel_row) AND ('0' & pixel_row <= cell_41y + cell_size)
				THEN
				CellDisplay(5, 0);
			ELSIF
				('0' & cell_42x <= pixel_column) AND ('0' & pixel_column <= cell_42x + cell_size) AND
				('0' & cell_42y <= pixel_row) AND ('0' & pixel_row <= cell_42y + cell_size)
				THEN
				CellDisplay(5, 1);
			ELSIF
				('0' & cell_43x <= pixel_column) AND ('0' & pixel_column <= cell_43x + cell_size) AND
				('0' & cell_43y <= pixel_row) AND ('0' & pixel_row <= cell_43y + cell_size)
				THEN
				CellDisplay(5, 2);
			ELSIF
				('0' & cell_44x <= pixel_column) AND ('0' & pixel_column <= cell_44x + cell_size) AND
				('0' & cell_44y <= pixel_row) AND ('0' & pixel_row <= cell_44y + cell_size)
				THEN
				CellDisplay(5, 3);
			ELSIF
				('0' & cell_45x <= pixel_column) AND ('0' & pixel_column <= cell_45x + cell_size) AND
				('0' & cell_45y <= pixel_row) AND ('0' & pixel_row <= cell_45y + cell_size)
				THEN
				CellDisplay(5, 4);
			ELSIF
				('0' & cell_46x <= pixel_column) AND ('0' & pixel_column <= cell_46x + cell_size) AND
				('0' & cell_46y <= pixel_row) AND ('0' & pixel_row <= cell_46y + cell_size)
				THEN
				CellDisplay(5, 5);
			ELSIF
				('0' & cell_47x <= pixel_column) AND ('0' & pixel_column <= cell_47x + cell_size) AND
				('0' & cell_47y <= pixel_row) AND ('0' & pixel_row <= cell_47y + cell_size)
				THEN
				CellDisplay(5, 6);
			ELSIF
				('0' & cell_48x <= pixel_column) AND ('0' & pixel_column <= cell_48x + cell_size) AND
				('0' & cell_48y <= pixel_row) AND ('0' & pixel_row <= cell_48y + cell_size)
				THEN
				CellDisplay(5, 7);
			ELSIF
				('0' & cell_49x <= pixel_column) AND ('0' & pixel_column <= cell_49x + cell_size) AND
				('0' & cell_49y <= pixel_row) AND ('0' & pixel_row <= cell_49y + cell_size)
				THEN
				CellDisplay(6, 0);
			ELSIF
				('0' & cell_50x <= pixel_column) AND ('0' & pixel_column <= cell_50x + cell_size) AND
				('0' & cell_50y <= pixel_row) AND ('0' & pixel_row <= cell_50y + cell_size)
				THEN
				CellDisplay(6, 1);
			ELSIF
				('0' & cell_51x <= pixel_column) AND ('0' & pixel_column <= cell_51x + cell_size) AND
				('0' & cell_51y <= pixel_row) AND ('0' & pixel_row <= cell_51y + cell_size)
				THEN
				CellDisplay(6, 2);
			ELSIF
				('0' & cell_52x <= pixel_column) AND ('0' & pixel_column <= cell_52x + cell_size) AND
				('0' & cell_52y <= pixel_row) AND ('0' & pixel_row <= cell_52y + cell_size)
				THEN
				CellDisplay(6, 3);
			ELSIF
				('0' & cell_53x <= pixel_column) AND ('0' & pixel_column <= cell_53x + cell_size) AND
				('0' & cell_53y <= pixel_row) AND ('0' & pixel_row <= cell_53y + cell_size)
				THEN
				CellDisplay(6, 4);
			ELSIF
				('0' & cell_54x <= pixel_column) AND ('0' & pixel_column <= cell_54x + cell_size) AND
				('0' & cell_54y <= pixel_row) AND ('0' & pixel_row <= cell_54y + cell_size)
				THEN
				CellDisplay(6, 5);
			ELSIF
				('0' & cell_55x <= pixel_column) AND ('0' & pixel_column <= cell_55x + cell_size) AND
				('0' & cell_55y <= pixel_row) AND ('0' & pixel_row <= cell_55y + cell_size)
				THEN
				CellDisplay(6, 6);
			ELSIF
				('0' & cell_56x <= pixel_column) AND ('0' & pixel_column <= cell_56x + cell_size) AND
				('0' & cell_56y <= pixel_row) AND ('0' & pixel_row <= cell_56y + cell_size)
				THEN
				CellDisplay(6, 7);
			ELSIF
				('0' & cell_57x <= pixel_column) AND ('0' & pixel_column <= cell_57x + cell_size) AND
				('0' & cell_57y <= pixel_row) AND ('0' & pixel_row <= cell_57y + cell_size)
				THEN
				CellDisplay(7, 0);
			ELSIF
				('0' & cell_58x <= pixel_column) AND ('0' & pixel_column <= cell_58x + cell_size) AND
				('0' & cell_58y <= pixel_row) AND ('0' & pixel_row <= cell_58y + cell_size)
				THEN
				CellDisplay(7, 1);
			ELSIF
				('0' & cell_59x <= pixel_column) AND ('0' & pixel_column <= cell_59x + cell_size) AND
				('0' & cell_59y <= pixel_row) AND ('0' & pixel_row <= cell_59y + cell_size)
				THEN
				CellDisplay(7, 2);
			ELSIF
				('0' & cell_60x <= pixel_column) AND ('0' & pixel_column <= cell_60x + cell_size) AND
				('0' & cell_60y <= pixel_row) AND ('0' & pixel_row <= cell_60y + cell_size)
				THEN
				CellDisplay(7, 3);
			ELSIF
				('0' & cell_61x <= pixel_column) AND ('0' & pixel_column <= cell_61x + cell_size) AND
				('0' & cell_61y <= pixel_row) AND ('0' & pixel_row <= cell_61y + cell_size)
				THEN
				CellDisplay(7, 4);
			ELSIF
				('0' & cell_62x <= pixel_column) AND ('0' & pixel_column <= cell_62x + cell_size) AND
				('0' & cell_62y <= pixel_row) AND ('0' & pixel_row <= cell_62y + cell_size)
				THEN
				CellDisplay(7, 5);
			ELSIF
				('0' & cell_63x <= pixel_column) AND ('0' & pixel_column <= cell_63x + cell_size) AND
				('0' & cell_63y <= pixel_row) AND ('0' & pixel_row <= cell_63y + cell_size)
				THEN
				CellDisplay(7, 6);
			ELSIF
				('0' & cell_64x <= pixel_column) AND ('0' & pixel_column <= cell_64x + cell_size) AND
				('0' & cell_64y <= pixel_row) AND ('0' & pixel_row <= cell_64y + cell_size)
				THEN
				CellDisplay(7, 7);
			ELSE
				Red <= grid_color(2);
				Green <= grid_color(1);
				Blue <= grid_color(0);
			END IF;
		END IF;
	END PROCESS RGB_Display;

END behavior;